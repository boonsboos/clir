module server

pub fn server() {
	
}