module server

import net

pub fn server() {
	
}