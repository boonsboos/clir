module main

import client
import util // imported so the settings work

fn main() {
	client.run()
}
