module main

import util

fn main() {

	if settings.server_mode {
		// server()
		println('server')
	} else {
		// client()
		println('client')
	}

}