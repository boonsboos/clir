module client

pub fn client() {
	
}